module testbench();
endmodule